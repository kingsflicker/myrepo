module test-file(input logic x, output log y)

  assign y = -x;

endmodule
